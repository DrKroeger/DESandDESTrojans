// The S MagicBoxes
module s_box(
input      [5:0] select_box0,
input      [5:0] select_box1,
input      [5:0] select_box2,
input      [5:0] select_box3,
input      [5:0] select_box4,
input      [5:0] select_box5,
input      [5:0] select_box6,
input      [5:0] select_box7,
output reg [3:0] s_out0,/* synthesis preserve */
output reg [3:0] s_out1,/* synthesis preserve */
output reg [3:0] s_out2,/* synthesis preserve */
output reg [3:0] s_out3,/* synthesis preserve */
output reg [3:0] s_out4,/* synthesis preserve */
output reg [3:0] s_out5,/* synthesis preserve */
output reg [3:0] s_out6,/* synthesis preserve */
output reg [3:0] s_out7 /* synthesis preserve */
);

always@(*) begin
case(select_box0)
//Box 0
  6'd0: s_out0 <= 4'hE;
  6'd1: s_out0 <= 4'h4;
  6'd2: s_out0 <= 4'hD;
  6'd3: s_out0 <= 4'h1;
  6'd4: s_out0 <= 4'h2;
  6'd5: s_out0 <= 4'hF;
  6'd6: s_out0 <= 4'hB;
  6'd7: s_out0 <= 4'h8;
  6'd8: s_out0 <= 4'h3;
  6'd9: s_out0 <= 4'hA;
  6'd10: s_out0 <= 4'h6;
  6'd11: s_out0 <= 4'hC;
  6'd12: s_out0 <= 4'h5;
  6'd13: s_out0 <= 4'h9;
  6'd14: s_out0 <= 4'h0;
  6'd15: s_out0 <= 4'h7;
  6'd16: s_out0 <= 4'h0;
  6'd17: s_out0 <= 4'hF;
  6'd18: s_out0 <= 4'h7;
  6'd19: s_out0 <= 4'h4;
  6'd20: s_out0 <= 4'hE;
  6'd21: s_out0 <= 4'h2;
  6'd22: s_out0 <= 4'hD;
  6'd23: s_out0 <= 4'h1;
  6'd24: s_out0 <= 4'hA;
  6'd25: s_out0 <= 4'h6;
  6'd26: s_out0 <= 4'hC;
  6'd27: s_out0 <= 4'hB;
  6'd28: s_out0 <= 4'h9;
  6'd29: s_out0 <= 4'h5;
  6'd30: s_out0 <= 4'h3;
  6'd31: s_out0 <= 4'h8;
  6'd32: s_out0 <= 4'h4;
  6'd33: s_out0 <= 4'h1;
  6'd34: s_out0 <= 4'hE;
  6'd35: s_out0 <= 4'h8;
  6'd36: s_out0 <= 4'hD;
  6'd37: s_out0 <= 4'h6;
  6'd38: s_out0 <= 4'h2;
  6'd39: s_out0 <= 4'hB;
  6'd40: s_out0 <= 4'hF;
  6'd41: s_out0 <= 4'hC;
  6'd42: s_out0 <= 4'h9;
  6'd43: s_out0 <= 4'h7;
  6'd44: s_out0 <= 4'h3;
  6'd45: s_out0 <= 4'hA;
  6'd46: s_out0 <= 4'h5;
  6'd47: s_out0 <= 4'h0;
  6'd48: s_out0 <= 4'hF;
  6'd49: s_out0 <= 4'hC;
  6'd50: s_out0 <= 4'h8;
  6'd51: s_out0 <= 4'h2;
  6'd52: s_out0 <= 4'h4;
  6'd53: s_out0 <= 4'h9;
  6'd54: s_out0 <= 4'h1;
  6'd55: s_out0 <= 4'h7;
  6'd56: s_out0 <= 4'h5;
  6'd57: s_out0 <= 4'hB;
  6'd58: s_out0 <= 4'h3;
  6'd59: s_out0 <= 4'hE;
  6'd60: s_out0 <= 4'hA;
  6'd61: s_out0 <= 4'h0;
  6'd62: s_out0 <= 4'h6;
  6'd63: s_out0 <= 4'hD;
  default: s_out0 <= 4'hX;
endcase

case(select_box1)
//Box 1
  6'd0: s_out1 <= 4'hF;
  6'd1: s_out1 <= 4'h1;
  6'd2: s_out1 <= 4'h8;
  6'd3: s_out1 <= 4'hE;
  6'd4: s_out1 <= 4'h6;
  6'd5: s_out1 <= 4'hB;
  6'd6: s_out1 <= 4'h3;
  6'd7: s_out1 <= 4'h4;
  6'd8: s_out1 <= 4'h9;
  6'd9: s_out1 <= 4'h7;
  6'd10: s_out1 <= 4'h2;
  6'd11: s_out1 <= 4'hD;
  6'd12: s_out1 <= 4'hC;
  6'd13: s_out1 <= 4'h0;
  6'd14: s_out1 <= 4'h5;
  6'd15: s_out1 <= 4'hA;
  6'd16: s_out1 <= 4'h3;
  6'd17: s_out1 <= 4'hD;
  6'd18: s_out1 <= 4'h4;
  6'd19: s_out1 <= 4'h7;
  6'd20: s_out1 <= 4'hF;
  6'd21: s_out1 <= 4'h2;
  6'd22: s_out1 <= 4'h8;
  6'd23: s_out1 <= 4'hE;
  6'd24: s_out1 <= 4'hC;
  6'd25: s_out1 <= 4'h0;
  6'd26: s_out1 <= 4'h1;
  6'd27: s_out1 <= 4'hA;
  6'd28: s_out1 <= 4'h6;
  6'd29: s_out1 <= 4'h9;
  6'd30: s_out1 <= 4'hB;
  6'd31: s_out1 <= 4'h5;
  6'd32: s_out1 <= 4'h0;
  6'd33: s_out1 <= 4'hE;
  6'd34: s_out1 <= 4'h7;
  6'd35: s_out1 <= 4'hB;
  6'd36: s_out1 <= 4'hA;
  6'd37: s_out1 <= 4'h4;
  6'd38: s_out1 <= 4'hD;
  6'd39: s_out1 <= 4'h1;
  6'd40: s_out1 <= 4'h5;
  6'd41: s_out1 <= 4'h8;
  6'd42: s_out1 <= 4'hC;
  6'd43: s_out1 <= 4'h6;
  6'd44: s_out1 <= 4'h9;
  6'd45: s_out1 <= 4'h3;
  6'd46: s_out1 <= 4'h2;
  6'd47: s_out1 <= 4'hF;
  6'd48: s_out1 <= 4'hD;
  6'd49: s_out1 <= 4'h8;
  6'd50: s_out1 <= 4'hA;
  6'd51: s_out1 <= 4'h1;
  6'd52: s_out1 <= 4'h3;
  6'd53: s_out1 <= 4'hF;
  6'd54: s_out1 <= 4'h4;
  6'd55: s_out1 <= 4'h2;
  6'd56: s_out1 <= 4'hB;
  6'd57: s_out1 <= 4'h6;
  6'd58: s_out1 <= 4'h7;
  6'd59: s_out1 <= 4'hC;
  6'd60: s_out1 <= 4'h0;
  6'd61: s_out1 <= 4'h5;
  6'd62: s_out1 <= 4'hE;
  6'd63: s_out1 <= 4'h9;
  default: s_out1 <= 4'hX;
endcase

case(select_box2)
//Box 2
  6'd0: s_out2 <= 4'hA;
  6'd1: s_out2 <= 4'h0;
  6'd2: s_out2 <= 4'h9;
  6'd3: s_out2 <= 4'hE;
  6'd4: s_out2 <= 4'h6;
  6'd5: s_out2 <= 4'h3;
  6'd6: s_out2 <= 4'hF;
  6'd7: s_out2 <= 4'h5;
  6'd8: s_out2 <= 4'h1;
  6'd9: s_out2 <= 4'hD;
  6'd10: s_out2 <= 4'hC;
  6'd11: s_out2 <= 4'h7;
  6'd12: s_out2 <= 4'hB;
  6'd13: s_out2 <= 4'h4;
  6'd14: s_out2 <= 4'h2;
  6'd15: s_out2 <= 4'h8;
  6'd16: s_out2 <= 4'hD;
  6'd17: s_out2 <= 4'h7;
  6'd18: s_out2 <= 4'h0;
  6'd19: s_out2 <= 4'h9;
  6'd20: s_out2 <= 4'h3;
  6'd21: s_out2 <= 4'h4;
  6'd22: s_out2 <= 4'h6;
  6'd23: s_out2 <= 4'hA;
  6'd24: s_out2 <= 4'h2;
  6'd25: s_out2 <= 4'h8;
  6'd26: s_out2 <= 4'h5;
  6'd27: s_out2 <= 4'hE;
  6'd28: s_out2 <= 4'hC;
  6'd29: s_out2 <= 4'hB;
  6'd30: s_out2 <= 4'hF;
  6'd31: s_out2 <= 4'h1;
  6'd32: s_out2 <= 4'hD;
  6'd33: s_out2 <= 4'h6;
  6'd34: s_out2 <= 4'h4;
  6'd35: s_out2 <= 4'h9;
  6'd36: s_out2 <= 4'h8;
  6'd37: s_out2 <= 4'hF;
  6'd38: s_out2 <= 4'h3;
  6'd39: s_out2 <= 4'h0;
  6'd40: s_out2 <= 4'hB;
  6'd41: s_out2 <= 4'h1;
  6'd42: s_out2 <= 4'h2;
  6'd43: s_out2 <= 4'hC;
  6'd44: s_out2 <= 4'h5;
  6'd45: s_out2 <= 4'hA;
  6'd46: s_out2 <= 4'hE;
  6'd47: s_out2 <= 4'h7;
  6'd48: s_out2 <= 4'h1;
  6'd49: s_out2 <= 4'hA;
  6'd50: s_out2 <= 4'hD;
  6'd51: s_out2 <= 4'h0;
  6'd52: s_out2 <= 4'h6;
  6'd53: s_out2 <= 4'h9;
  6'd54: s_out2 <= 4'h8;
  6'd55: s_out2 <= 4'h7;
  6'd56: s_out2 <= 4'h4;
  6'd57: s_out2 <= 4'hF;
  6'd58: s_out2 <= 4'hE;
  6'd59: s_out2 <= 4'h3;
  6'd60: s_out2 <= 4'hB;
  6'd61: s_out2 <= 4'h5;
  6'd62: s_out2 <= 4'h2;
  6'd63: s_out2 <= 4'hC;
  default: s_out2 <= 4'hX;
endcase

case(select_box3)
//Box 3
  6'd0: s_out3 <= 4'h7;
  6'd1: s_out3 <= 4'hD;
  6'd2: s_out3 <= 4'hE;
  6'd3: s_out3 <= 4'h3;
  6'd4: s_out3 <= 4'h0;
  6'd5: s_out3 <= 4'h6;
  6'd6: s_out3 <= 4'h9;
  6'd7: s_out3 <= 4'hA;
  6'd8: s_out3 <= 4'h1;
  6'd9: s_out3 <= 4'h2;
  6'd10: s_out3 <= 4'h8;
  6'd11: s_out3 <= 4'h5;
  6'd12: s_out3 <= 4'hB;
  6'd13: s_out3 <= 4'hC;
  6'd14: s_out3 <= 4'h4;
  6'd15: s_out3 <= 4'hF;
  6'd16: s_out3 <= 4'hD;
  6'd17: s_out3 <= 4'h8;
  6'd18: s_out3 <= 4'hB;
  6'd19: s_out3 <= 4'h5;
  6'd20: s_out3 <= 4'h6;
  6'd21: s_out3 <= 4'hF;
  6'd22: s_out3 <= 4'h0;
  6'd23: s_out3 <= 4'h3;
  6'd24: s_out3 <= 4'h4;
  6'd25: s_out3 <= 4'h7;
  6'd26: s_out3 <= 4'h2;
  6'd27: s_out3 <= 4'hC;
  6'd28: s_out3 <= 4'h1;
  6'd29: s_out3 <= 4'hA;
  6'd30: s_out3 <= 4'hE;
  6'd31: s_out3 <= 4'h9;
  6'd32: s_out3 <= 4'hA;
  6'd33: s_out3 <= 4'h6;
  6'd34: s_out3 <= 4'h9;
  6'd35: s_out3 <= 4'h0;
  6'd36: s_out3 <= 4'hC;
  6'd37: s_out3 <= 4'hB;
  6'd38: s_out3 <= 4'h7;
  6'd39: s_out3 <= 4'hD;
  6'd40: s_out3 <= 4'hF;
  6'd41: s_out3 <= 4'h1;
  6'd42: s_out3 <= 4'h3;
  6'd43: s_out3 <= 4'hE;
  6'd44: s_out3 <= 4'h5;
  6'd45: s_out3 <= 4'h2;
  6'd46: s_out3 <= 4'h8;
  6'd47: s_out3 <= 4'h4;
  6'd48: s_out3 <= 4'h3;
  6'd49: s_out3 <= 4'hF;
  6'd50: s_out3 <= 4'h0;
  6'd51: s_out3 <= 4'h6;
  6'd52: s_out3 <= 4'hA;
  6'd53: s_out3 <= 4'h1;
  6'd54: s_out3 <= 4'hD;
  6'd55: s_out3 <= 4'h8;
  6'd56: s_out3 <= 4'h9;
  6'd57: s_out3 <= 4'h4;
  6'd58: s_out3 <= 4'h5;
  6'd59: s_out3 <= 4'hB;
  6'd60: s_out3 <= 4'hC;
  6'd61: s_out3 <= 4'h7;
  6'd62: s_out3 <= 4'h2;
  6'd63: s_out3 <= 4'hE;
  default: s_out3 <= 4'hX;
endcase

case(select_box4)
//Box 4
  6'd0: s_out4 <= 4'h2;
  6'd1: s_out4 <= 4'hC;
  6'd2: s_out4 <= 4'h4;
  6'd3: s_out4 <= 4'h1;
  6'd4: s_out4 <= 4'h7;
  6'd5: s_out4 <= 4'hA;
  6'd6: s_out4 <= 4'hB;
  6'd7: s_out4 <= 4'h6;
  6'd8: s_out4 <= 4'h8;
  6'd9: s_out4 <= 4'h5;
  6'd10: s_out4 <= 4'h3;
  6'd11: s_out4 <= 4'hF;
  6'd12: s_out4 <= 4'hD;
  6'd13: s_out4 <= 4'h0;
  6'd14: s_out4 <= 4'hE;
  6'd15: s_out4 <= 4'h9;
  6'd16: s_out4 <= 4'hE;
  6'd17: s_out4 <= 4'hB;
  6'd18: s_out4 <= 4'h2;
  6'd19: s_out4 <= 4'hC;
  6'd20: s_out4 <= 4'h4;
  6'd21: s_out4 <= 4'h7;
  6'd22: s_out4 <= 4'hD;
  6'd23: s_out4 <= 4'h1;
  6'd24: s_out4 <= 4'h5;
  6'd25: s_out4 <= 4'h0;
  6'd26: s_out4 <= 4'hF;
  6'd27: s_out4 <= 4'hA;
  6'd28: s_out4 <= 4'h3;
  6'd29: s_out4 <= 4'h9;
  6'd30: s_out4 <= 4'h8;
  6'd31: s_out4 <= 4'h6;
  6'd32: s_out4 <= 4'h4;
  6'd33: s_out4 <= 4'h2;
  6'd34: s_out4 <= 4'h1;
  6'd35: s_out4 <= 4'hB;
  6'd36: s_out4 <= 4'hA;
  6'd37: s_out4 <= 4'hD;
  6'd38: s_out4 <= 4'h7;
  6'd39: s_out4 <= 4'h8;
  6'd40: s_out4 <= 4'hF;
  6'd41: s_out4 <= 4'h9;
  6'd42: s_out4 <= 4'hC;
  6'd43: s_out4 <= 4'h5;
  6'd44: s_out4 <= 4'h6;
  6'd45: s_out4 <= 4'h3;
  6'd46: s_out4 <= 4'h0;
  6'd47: s_out4 <= 4'hE;
  6'd48: s_out4 <= 4'hB;
  6'd49: s_out4 <= 4'h8;
  6'd50: s_out4 <= 4'hC;
  6'd51: s_out4 <= 4'h7;
  6'd52: s_out4 <= 4'h1;
  6'd53: s_out4 <= 4'hE;
  6'd54: s_out4 <= 4'h2;
  6'd55: s_out4 <= 4'hD;
  6'd56: s_out4 <= 4'h6;
  6'd57: s_out4 <= 4'hF;
  6'd58: s_out4 <= 4'h0;
  6'd59: s_out4 <= 4'h9;
  6'd60: s_out4 <= 4'hA;
  6'd61: s_out4 <= 4'h4;
  6'd62: s_out4 <= 4'h5;
  6'd63: s_out4 <= 4'h3;
  default: s_out4 <= 4'hX;
endcase

case(select_box5)
//Box 5
  6'd0: s_out5 <= 4'hC;
  6'd1: s_out5 <= 4'h1;
  6'd2: s_out5 <= 4'hA;
  6'd3: s_out5 <= 4'hF;
  6'd4: s_out5 <= 4'h9;
  6'd5: s_out5 <= 4'h2;
  6'd6: s_out5 <= 4'h6;
  6'd7: s_out5 <= 4'h8;
  6'd8: s_out5 <= 4'h0;
  6'd9: s_out5 <= 4'hD;
  6'd10: s_out5 <= 4'h3;
  6'd11: s_out5 <= 4'h4;
  6'd12: s_out5 <= 4'hE;
  6'd13: s_out5 <= 4'h7;
  6'd14: s_out5 <= 4'h5;
  6'd15: s_out5 <= 4'hB;
  6'd16: s_out5 <= 4'hA;
  6'd17: s_out5 <= 4'hF;
  6'd18: s_out5 <= 4'h4;
  6'd19: s_out5 <= 4'h2;
  6'd20: s_out5 <= 4'h7;
  6'd21: s_out5 <= 4'hC;
  6'd22: s_out5 <= 4'h9;
  6'd23: s_out5 <= 4'h5;
  6'd24: s_out5 <= 4'h6;
  6'd25: s_out5 <= 4'h1;
  6'd26: s_out5 <= 4'hD;
  6'd27: s_out5 <= 4'hE;
  6'd28: s_out5 <= 4'h0;
  6'd29: s_out5 <= 4'hB;
  6'd30: s_out5 <= 4'h3;
  6'd31: s_out5 <= 4'h8;
  6'd32: s_out5 <= 4'h9;
  6'd33: s_out5 <= 4'hE;
  6'd34: s_out5 <= 4'hF;
  6'd35: s_out5 <= 4'h5;
  6'd36: s_out5 <= 4'h2;
  6'd37: s_out5 <= 4'h8;
  6'd38: s_out5 <= 4'hC;
  6'd39: s_out5 <= 4'h3;
  6'd40: s_out5 <= 4'h7;
  6'd41: s_out5 <= 4'h0;
  6'd42: s_out5 <= 4'h4;
  6'd43: s_out5 <= 4'hA;
  6'd44: s_out5 <= 4'h1;
  6'd45: s_out5 <= 4'hD;
  6'd46: s_out5 <= 4'hB;
  6'd47: s_out5 <= 4'h6;
  6'd48: s_out5 <= 4'h4;
  6'd49: s_out5 <= 4'h3;
  6'd50: s_out5 <= 4'h2;
  6'd51: s_out5 <= 4'hC;
  6'd52: s_out5 <= 4'h9;
  6'd53: s_out5 <= 4'h5;
  6'd54: s_out5 <= 4'hF;
  6'd55: s_out5 <= 4'hA;
  6'd56: s_out5 <= 4'hB;
  6'd57: s_out5 <= 4'hE;
  6'd58: s_out5 <= 4'h1;
  6'd59: s_out5 <= 4'h7;
  6'd60: s_out5 <= 4'h6;
  6'd61: s_out5 <= 4'h0;
  6'd62: s_out5 <= 4'h8;
  6'd63: s_out5 <= 4'hD;
  default: s_out5 <= 4'hX;
endcase

case(select_box6)
//Box 6
  6'd0: s_out6 <= 4'h4;
  6'd1: s_out6 <= 4'hB;
  6'd2: s_out6 <= 4'h2;
  6'd3: s_out6 <= 4'hE;
  6'd4: s_out6 <= 4'hF;
  6'd5: s_out6 <= 4'h0;
  6'd6: s_out6 <= 4'h8;
  6'd7: s_out6 <= 4'hD;
  6'd8: s_out6 <= 4'h3;
  6'd9: s_out6 <= 4'hC;
  6'd10: s_out6 <= 4'h9;
  6'd11: s_out6 <= 4'h7;
  6'd12: s_out6 <= 4'h5;
  6'd13: s_out6 <= 4'hA;
  6'd14: s_out6 <= 4'h6;
  6'd15: s_out6 <= 4'h1;
  6'd16: s_out6 <= 4'hD;
  6'd17: s_out6 <= 4'h0;
  6'd18: s_out6 <= 4'hB;
  6'd19: s_out6 <= 4'h7;
  6'd20: s_out6 <= 4'h4;
  6'd21: s_out6 <= 4'h9;
  6'd22: s_out6 <= 4'h1;
  6'd23: s_out6 <= 4'hA;
  6'd24: s_out6 <= 4'hE;
  6'd25: s_out6 <= 4'h3;
  6'd26: s_out6 <= 4'h5;
  6'd27: s_out6 <= 4'hC;
  6'd28: s_out6 <= 4'h2;
  6'd29: s_out6 <= 4'hF;
  6'd30: s_out6 <= 4'h8;
  6'd31: s_out6 <= 4'h6;
  6'd32: s_out6 <= 4'h1;
  6'd33: s_out6 <= 4'h4;
  6'd34: s_out6 <= 4'hB;
  6'd35: s_out6 <= 4'hD;
  6'd36: s_out6 <= 4'hC;
  6'd37: s_out6 <= 4'h3;
  6'd38: s_out6 <= 4'h7;
  6'd39: s_out6 <= 4'hE;
  6'd40: s_out6 <= 4'hA;
  6'd41: s_out6 <= 4'hF;
  6'd42: s_out6 <= 4'h6;
  6'd43: s_out6 <= 4'h8;
  6'd44: s_out6 <= 4'h0;
  6'd45: s_out6 <= 4'h5;
  6'd46: s_out6 <= 4'h9;
  6'd47: s_out6 <= 4'h2;
  6'd48: s_out6 <= 4'h6;
  6'd49: s_out6 <= 4'hB;
  6'd50: s_out6 <= 4'hD;
  6'd51: s_out6 <= 4'h8;
  6'd52: s_out6 <= 4'h1;
  6'd53: s_out6 <= 4'h4;
  6'd54: s_out6 <= 4'hA;
  6'd55: s_out6 <= 4'h7;
  6'd56: s_out6 <= 4'h9;
  6'd57: s_out6 <= 4'h5;
  6'd58: s_out6 <= 4'h0;
  6'd59: s_out6 <= 4'hF;
  6'd60: s_out6 <= 4'hE;
  6'd61: s_out6 <= 4'h2;
  6'd62: s_out6 <= 4'h3;
  6'd63: s_out6 <= 4'hC;
  default: s_out6 <= 4'hX;
endcase

case(select_box7)
//Box 7
  6'd0: s_out7 <= 4'hD;
  6'd1: s_out7 <= 4'h2;
  6'd2: s_out7 <= 4'h8;
  6'd3: s_out7 <= 4'h4;
  6'd4: s_out7 <= 4'h6;
  6'd5: s_out7 <= 4'hF;
  6'd6: s_out7 <= 4'hB;
  6'd7: s_out7 <= 4'h1;
  6'd8: s_out7 <= 4'hA;
  6'd9: s_out7 <= 4'h9;
  6'd10: s_out7 <= 4'h3;
  6'd11: s_out7 <= 4'hE;
  6'd12: s_out7 <= 4'h5;
  6'd13: s_out7 <= 4'h0;
  6'd14: s_out7 <= 4'hC;
  6'd15: s_out7 <= 4'h7;
  6'd16: s_out7 <= 4'h1;
  6'd17: s_out7 <= 4'hF;
  6'd18: s_out7 <= 4'hD;
  6'd19: s_out7 <= 4'h8;
  6'd20: s_out7 <= 4'hA;
  6'd21: s_out7 <= 4'h3;
  6'd22: s_out7 <= 4'h7;
  6'd23: s_out7 <= 4'h4;
  6'd24: s_out7 <= 4'hC;
  6'd25: s_out7 <= 4'h5;
  6'd26: s_out7 <= 4'h6;
  6'd27: s_out7 <= 4'hB;
  6'd28: s_out7 <= 4'h0;
  6'd29: s_out7 <= 4'hE;
  6'd30: s_out7 <= 4'h9;
  6'd31: s_out7 <= 4'h2;
  6'd32: s_out7 <= 4'h7;
  6'd33: s_out7 <= 4'hB;
  6'd34: s_out7 <= 4'h4;
  6'd35: s_out7 <= 4'h1;
  6'd36: s_out7 <= 4'h9;
  6'd37: s_out7 <= 4'hC;
  6'd38: s_out7 <= 4'hE;
  6'd39: s_out7 <= 4'h2;
  6'd40: s_out7 <= 4'h0;
  6'd41: s_out7 <= 4'h6;
  6'd42: s_out7 <= 4'hA;
  6'd43: s_out7 <= 4'hD;
  6'd44: s_out7 <= 4'hF;
  6'd45: s_out7 <= 4'h3;
  6'd46: s_out7 <= 4'h5;
  6'd47: s_out7 <= 4'h8;
  6'd48: s_out7 <= 4'h2;
  6'd49: s_out7 <= 4'h1;
  6'd50: s_out7 <= 4'hE;
  6'd51: s_out7 <= 4'h7;
  6'd52: s_out7 <= 4'h4;
  6'd53: s_out7 <= 4'hA;
  6'd54: s_out7 <= 4'h8;
  6'd55: s_out7 <= 4'hD;
  6'd56: s_out7 <= 4'hF;
  6'd57: s_out7 <= 4'hC;
  6'd58: s_out7 <= 4'h9;
  6'd59: s_out7 <= 4'h0;
  6'd60: s_out7 <= 4'h3;
  6'd61: s_out7 <= 4'h5;
  6'd62: s_out7 <= 4'h6;
  6'd63: s_out7 <= 4'hB;
  default: s_out7 <= 4'hX;
endcase

end
 
endmodule
